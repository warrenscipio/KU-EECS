`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    09:21:39 03/14/2013 
// Design Name: 
// Module Name:    twobitxor 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module twobitxor(A, B, C, F);
    input [0:0] A;
    input [0:0] B;
    input [0:0] C;
    output [0:0] F;


endmodule
