----------------------------------------------------------------------------------
-- Company: 
-- Engineer: Warren Scipio
-- 
-- Create Date:    09:50:16 03/07/2013 
-- Design Name: 
-- Module Name:    toplevel(hard) - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity toplevel(hard) is


end toplevel(hard);

architecture Behavioral of toplevel(hard) is

begin


end Behavioral;

